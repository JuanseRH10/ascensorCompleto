library verilog;
use verilog.vl_types.all;
entity capturarLlego_vlg_vec_tst is
end capturarLlego_vlg_vec_tst;
