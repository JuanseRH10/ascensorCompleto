library verilog;
use verilog.vl_types.all;
entity alarmas_vlg_vec_tst is
end alarmas_vlg_vec_tst;
