library verilog;
use verilog.vl_types.all;
entity registrosBotones_vlg_vec_tst is
end registrosBotones_vlg_vec_tst;
