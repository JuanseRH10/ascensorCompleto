library verilog;
use verilog.vl_types.all;
entity detectorPiso_vlg_vec_tst is
end detectorPiso_vlg_vec_tst;
