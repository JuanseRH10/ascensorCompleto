library verilog;
use verilog.vl_types.all;
entity controlPuerta_vlg_vec_tst is
end controlPuerta_vlg_vec_tst;
