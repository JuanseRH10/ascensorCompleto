library verilog;
use verilog.vl_types.all;
entity detectorBoton_vlg_vec_tst is
end detectorBoton_vlg_vec_tst;
