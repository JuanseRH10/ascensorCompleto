library verilog;
use verilog.vl_types.all;
entity actualizarPiso_vlg_vec_tst is
end actualizarPiso_vlg_vec_tst;
