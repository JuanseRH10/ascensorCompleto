library verilog;
use verilog.vl_types.all;
entity div_frec_vlg_vec_tst is
end div_frec_vlg_vec_tst;
