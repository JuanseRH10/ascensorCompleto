library verilog;
use verilog.vl_types.all;
entity controlContadores_vlg_vec_tst is
end controlContadores_vlg_vec_tst;
