library verilog;
use verilog.vl_types.all;
entity contadorPersonas_vlg_vec_tst is
end contadorPersonas_vlg_vec_tst;
