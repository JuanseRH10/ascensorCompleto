library verilog;
use verilog.vl_types.all;
entity contadorSeg_vlg_vec_tst is
end contadorSeg_vlg_vec_tst;
