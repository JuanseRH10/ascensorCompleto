library verilog;
use verilog.vl_types.all;
entity detectorCambio_vlg_vec_tst is
end detectorCambio_vlg_vec_tst;
