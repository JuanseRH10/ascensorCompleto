library verilog;
use verilog.vl_types.all;
entity movimientoAscensor_vlg_vec_tst is
end movimientoAscensor_vlg_vec_tst;
