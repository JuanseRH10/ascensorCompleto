library verilog;
use verilog.vl_types.all;
entity comparadorNbits_vlg_vec_tst is
end comparadorNbits_vlg_vec_tst;
