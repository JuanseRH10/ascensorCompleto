library verilog;
use verilog.vl_types.all;
entity decun_vlg_vec_tst is
end decun_vlg_vec_tst;
