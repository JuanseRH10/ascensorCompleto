library verilog;
use verilog.vl_types.all;
entity contadorGenerico_vlg_vec_tst is
end contadorGenerico_vlg_vec_tst;
