library verilog;
use verilog.vl_types.all;
entity capturarLlego_vlg_check_tst is
    port(
        llego_capturado : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end capturarLlego_vlg_check_tst;
