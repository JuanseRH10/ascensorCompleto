library verilog;
use verilog.vl_types.all;
entity comparadorNbits_vlg_check_tst is
    port(
        AiguB           : in     vl_logic;
        AmayB           : in     vl_logic;
        AmenB           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end comparadorNbits_vlg_check_tst;
