library verilog;
use verilog.vl_types.all;
entity sensorPersonas_vlg_vec_tst is
end sensorPersonas_vlg_vec_tst;
