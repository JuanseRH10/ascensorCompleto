library verilog;
use verilog.vl_types.all;
entity controlAscensor_vlg_vec_tst is
end controlAscensor_vlg_vec_tst;
