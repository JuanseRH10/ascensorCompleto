library verilog;
use verilog.vl_types.all;
entity div_frec_vlg_check_tst is
    port(
        out1            : in     vl_logic;
        out2            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end div_frec_vlg_check_tst;
