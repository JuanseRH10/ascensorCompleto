library verilog;
use verilog.vl_types.all;
entity detectorCambio_vlg_check_tst is
    port(
        salida          : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end detectorCambio_vlg_check_tst;
